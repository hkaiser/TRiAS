���Z     @  4   I�         &                                       B
    �                                                     !   �   �� 	   ,          � Project@Options� -�   !�     7   \+ 	   -          � File@@Version2.1  � 1.1     (                                                          �   f   TOPIC VERSION OBJARRAY BROWSE_SEQUENCE BUILD_TAG CONTEX    link viewHandles 7                                            _ISECT_iterator _AE_Sorter _AE_mark _SysInfoFlags _outside_   Metafile VbPicture VbVarArray VeRec ViewEngine WinImage _AE   r VB_Historian VB_View VbCurrency VbDibBitmap VbFixArray Vb	   ng SystemDatabase TextFileDatabase TrashCollector TreeWalke
   Real RecordMark RuleSpecifier SchemaEngine SmartString Stri   adStream NamedData NamedMonad NilMonad Number Presentation    Dictionary Integer LogStream Monad MonadArray MonadFile Mon   tion Bcd36 Boolean ClassDesc ClassMethod ComboElement Date    Set AdRec AeAccessSet AgilityDatabase ArrayDatabase Associa   ]  YAccessCombo AccessEngine AccessItem AccessRule Access                    .       ,       )       #       �       �       &�       (      @)      E      Q�       uP      y      |}      ~�      ��      �*      �v      ��      ��      û      ��      �      �       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  n0    !� BuildAll!� 2!� Inhaltsverzeichnis!�% Copyright � 1991    Title , Arial ,  18 ,  180 ,  250 ,  40 ,  40 ,  0 , -1 , "   ['  �� 	   ,          � F1ProjectStyle2-'-�  � !�F�   92), 0!�3 "Index", ( 509, 0, 509, 1020), , , (192,192,192),$   2,192), 0!�4 "Glossary", ( 0, 0, 506, 1017), , , (192,192,1%   , (192,192,192), 0!�. "", ( 0, 505, 1018, 505), , , (192,19&   4, 453), , , (192,192,192), 0!�, "", ( 0, 0, 1018, 505), , '   $ "TRiAS� FAQ", , , , (192,192,192), 0!�. "", ( 471, 29, 51(   d  �u 	   -          � F1ProjectWindows5-�   !�    �  !�  !�  !�  !�  !�  !�                                  *     !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !+   �   � 	   -          � F1ProjectButtons^ -�   !�  �� aktiviertes Objekt,(Global), 2,Ein Objekt, welches nach -   �  �� 	   .          � F1ProjectGlossary�-�  6 !�    No!�  !�
 TRiAS� FAQ!� 1!�  !�  !�  !�                  /   5 uve GmbH FEZ Potsdam!�  !�  !�  !� 0!�  !�  !� 0!� 0!�@    0 , None , !�F Title , Arial ,  18 ,  120 ,  250 ,  40 ,  A   ,  180 ,  250 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�H Headi2   60 ,  20 ,  0 , -1 ,  0 , None , !�H Heading , Arial ,  12 3   1 ,  0 , None , !�H Heading , Arial ,  12 ,  180 ,  250 ,  4   �H Heading , Arial ,  12 ,  180 ,  250 ,  60 ,  20 ,  0 , -5   l ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !6   50 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�J Paragraph , Aria7   0 ,  0 ,  0 , Box , !�J Paragraph , Arial ,  10 ,  180 ,  28    ����Paragraph2 , Arial ,  10 ,  600 ,  250 ,  20 ,  60 ,  9   ,  10 ,  400 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�N:   0 ,  60 ,  0 ,  0 ,  0 , None , !�O ����Paragraph1 , Arial ;     0 , None , !�J Paragraph , Arial ,  10 ,  180 ,  250 ,  2<   F Title , Arial ,  18 ,  120 ,  250 ,  40 ,  40 ,  0 , -1 ,=    ,  18 ,  120 ,  250 ,  40 ,  40 ,  0 , -1 ,  0 , None , !�>     250 ,  40 ,  40 ,  0 , -1 ,  0 , None , !�F Title , Arial?   40 ,  0 , -1 ,  0 , None , !�F Title , Arial ,  18 ,  120 ,P   ng , Arial ,  12 ,  180 ,  250 ,  60 ,  20 ,  0 , -1 ,  0 ,Q   Arial ,  10 ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 ,  0 , NonB    250 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�L Jump Label , C   0 ,  0 ,  0 , None , !�L Jump Label , Arial ,  10 ,  180 , D   !�L Jump Label , Arial ,  10 ,  180 ,  250 ,  20 ,  20 ,  1E   l ,  10 ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 ,  0 , None , F    ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�L Jump Label , AriaG   -1 , -1 , None , !�L Jump Label , Arial ,  10 ,  180 ,  250H   Sub Heading , Arial ,  12 ,  180 ,  250 ,  40 ,  20 ,  0 , I     12 ,  180 ,  250 ,  40 ,  20 ,  0 , -1 , -1 , None , !�L J    40 ,  20 ,  0 , -1 , -1 , None , !�L Sub Heading , Arial ,K    -1 , None , !�L Sub Heading , Arial ,  12 ,  180 ,  250 , L   eading1 , Arial ,  12 ,  180 ,  250 ,  40 ,  20 ,  1 , -1 ,M   80 ,  250 ,  40 ,  20 ,  0 , -1 , -1 , None , !�Q ����Sub HN    ,  0 , -1 ,  0 , None , !�L Sub Heading , Arial ,  12 ,  1O    None , !�H Heading , Arial ,  12 ,  180 ,  250 ,  60 ,  20`   e , !�N Mono Spaced , Courier ,  10 ,  180 ,  250 ,  20 ,  a   tmap Paragraph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0R   10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�Q BiS   60 ,  0 ,  0 ,  0 , None , !�Q Bitmap Paragraph , Arial ,  T    , None , !�H Footnote , Arial ,  8 ,  180 ,  250 ,  20 ,  U   tnote , Arial ,  8 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0V   8 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�H FooW     20 ,  60 ,  0 ,  0 ,  0 , None , !�H Footnote , Arial ,  X     0 ,  0 , None , !�H Footnote , Arial ,  8 ,  180 ,  250 ,Y    !�H Footnote , Arial ,  8 ,  180 ,  250 ,  20 ,  60 ,  0 ,Z   ier ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None ,[    ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�N Mono Spaced , Cour\   ,  0 , None , !�N Mono Spaced , Courier ,  10 ,  180 ,  250]   Spaced , Courier ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ^   ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�N Mono _   60 ,  0 ,  0 ,  0 , None , !�N Mono Spaced , Courier ,  10 p    ,  0 ,  0 , None , !�Q Bitmap Paragraph , Arial ,  10 ,  1q   ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�G Bulleb    20 ,  60 ,  0 ,  0 , -1 , None , !�G Bullet , Arial ,  10 c     0 , None , !�L ����Bullet1 , Arial ,  10 ,  180 ,  250 , d    Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,e   ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�Gf     60 ,  0 ,  0 ,  0 , None , !�R Bitmap Jump Label , Arial g   , !�R Bitmap Jump Label , Arial ,  10 ,  180 ,  250 ,  20 ,h   rial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None i    20 ,  60 ,  0 ,  0 ,  0 , None , !�R Bitmap Jump Label , Aj   None , !�R Bitmap Jump Label , Arial ,  10 ,  180 ,  250 , k   l , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , l   50 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Bitmap Jump Labem     0 , None , !�Q Bitmap Paragraph , Arial ,  10 ,  180 ,  2n   ragraph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,o   80 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�Q Bitmap Pa��   t , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , �    , None , !�M Outline Node , Arial ,  10 ,  180 ,  250 ,  2r   Node , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0s   180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�M Outline t    ,  0 ,  0 ,  0 , None , !�M Outline Node , Arial ,  10 ,  u    , !�M Outline Node , Arial ,  10 ,  180 ,  250 ,  20 ,  60v   Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , Nonew   250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�M Outline Node , x     0 , None , !�R Enumerated Bullet , Arial ,  10 ,  180 ,  y    Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,z   0 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Enumerated{     0 ,  0 , None , !�R Enumerated Bullet , Arial ,  10 ,  18|   rated Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,}   ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Enume~     0 ,  0 ,  0 , None , !�R Enumerated Bullet , Arial ,  10    None , !�G Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,�   0 ,  60 ,  0 ,  0 ,  0 , None , !�M Outline Leaf , Arial , �   e , !�S Index Letter Label , Arial ,  12 ,  180 ,  250 ,  2�    Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , Non�     20 ,  60 ,  0 ,  0 ,  0 , None , !�S Index Letter Label ,�   0 ,  0 ,  0 , None , !�E Line , Arial ,  10 ,  180 ,  250 ,�   None , !�E Line , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  �   e , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , �   0 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�E Lin�   0 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�E Line , Arial ,  1�   ,  0 ,  0 ,  0 , None , !�E Line , Arial ,  10 ,  180 ,  25�   , !�M Outline Leaf , Arial ,  10 ,  180 ,  250 ,  20 ,  60 �   rial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None �   50 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�M Outline Leaf , A�    0 ,  0 , None , !�M Outline Leaf , Arial ,  10 ,  180 ,  2�   utline Leaf , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 , �    10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�M O�   0 ,  60 ,  0 , -1 ,  0 , None , !�S Index Letter Label , Ar�    180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�V Glossar�   -1 ,  0 , None , !�V Glossary Letter Label , Arial ,  12 , �   etter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , �   0 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�V Glossary L�   ,  0 , None , !�V Glossary Letter Label , Arial ,  12 ,  18�   �F Index , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 �   l ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�   ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Index , Aria�    60 ,  0 ,  0 ,  0 , None , !�F Index , Arial ,  10 ,  180 �     0 , None , !�F Index , Arial ,  10 ,  180 ,  250 ,  20 , �   F Index , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,�    ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !��     60 ,  0 , -1 ,  0 , None , !�S Index Letter Label , Arial�    !�S Index Letter Label , Arial ,  12 ,  180 ,  250 ,  20 ,�   ial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None ,B�   y Letter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0�   50 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�D Bar , Arial ,  1�   ,  0 ,  0 ,  0 , None , !�F Image , Arial ,  10 ,  180 ,  2�   , None , !�F Image , Arial ,  10 ,  180 ,  250 ,  20 ,  60 �   age , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 �   10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Im�   0 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Image , Arial ,  �     0 ,  0 ,  0 , None , !�F Image , Arial ,  10 ,  180 ,  25�   ne , !�I Glossary , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,�   , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , No�   80 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�I Glossary �    60 ,  0 ,  0 ,  0 , None , !�I Glossary , Arial ,  10 ,  1�    , None , !�I Glossary , Arial ,  10 ,  180 ,  250 ,  20 , �   sary , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0�    ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�I Glos�    , -1 ,  0 , None , !�V Glossary Letter Label , Arial ,  12�   0 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�D Bar�   ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,�   1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  �    Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !��   al ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�;  ,�     10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�;  , Ari�   ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,�   1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  �    Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !��   al ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�;  ,�     10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�;  , Ari�   0 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�;  , Arial ,�   0 ,  60 ,  0 ,  0 ,  0 , None , !�D Bar , Arial ,  10 ,  18�   ,  0 ,  0 , None , !�D Bar , Arial ,  10 ,  180 ,  250 ,  2�   one , !�D Bar , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 �    , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , Nn�     10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�;  , Ari�     10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�;  , Ari�   ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,�   1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  �    Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !��   al ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�;  ,�     10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�;  , Ari�   ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,�   1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  �    Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !��   al ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�;  ,�     10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�;  , Ari�   ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,�   1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  �    Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !��   al ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�;  ,�   al ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�;  ,�   �   M��� 
&  + 2 G     � Topic@Anhang A  �    � �     L��� 
(  7 > S     � Topic@Stichwortverzeichnis     /Style /Just L!� /X /Style /Just L  
q �  � 1004     �     �  �� 	\�   N -�   !� /T N /Just L /Text Index!� /Z N�   � �     �  ��6S     �  �� =h   
  � Index�� Lx   �   �   ��� 
  ( / D     � Topic@Index  �    �  �    L!� /Y /Style /Just L  
� �  � 1014                   �    N /Just L /Text Stichwortverzeichnis!� /Z N /Style /Just     T_STRING HELP_MACRO KEYWORDS TOPIC_TITLE NOTE              �   tichwortverzeichnis�� [�     �  �� 	k�   ] -�   !�' /T�     �    �  ��     �  ��Eb     �  �� L�     � Sk    10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�;  , Ari�   ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,�   1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  �    Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !���    �� �     �  ��9V     �  �� @n     � Anhang A�� �   e und Identifikator vor. Begrifflich sind beide entsprechen�   S� eine faktische inhaltlice Gleichstellung von Objektklass�   tklassen ist der Identifikator. Zur Zeit findet man in TRiA�   wendete Kriterium der Zusammenfassung von Objekten zu Objek�   ktklassen�� X�     �  �� 	h�  -�   !�  /T N /Just L4   /Text Objektklassen!� /P /Just L /Text !�k /L /Jump Was i�    Linienobjekt!� /B /Just L /Text Fl�chenobjekt!� /B /Just     � 1001                                                      L /Text Textobjekt!�� /P /Just L /Text Ein Objekt bietet d�     �  	  � 1011   �  ��>_     �  �� I|     � Obje�   �  �x�� 
u  0 7 P     � Topic@Objektklassen  �  �   schen oder anderen Kriterien.����Das wohl am h�ufigsten ver�   ammenfassung beliebiger Objekte nach geometrischen, themati�   A!�, /P /Just L /Text Insert Appendix A text here  
w � �   O~     �  �� 	_�   U -�   !� /T N /Just L /Text Anhang 8  d ihrem Sinn verwendet.����Die Objektklasse eines Objektes      0!�                                                          �    �  	  � 1016   �  ��C�   A  �< Raumbezug;Texto                                                               �   popup Main /Just L /Text Darstellung von Objekten (Farbe, S�   ignaturen etc.)!�Z /L /Jump Doppelte Menupunkte /Link /Macr�   o /Play /popup /Just L /Text Doppelte Menupunkte ?!�c /L /J�   ump Komandozeilenparameter /Link /Macro /Play /popup Main /�   Just L /Text Komandozeilenparameter!�[ /L /Jump Koordinaten�   systeme /Link /Macro /Play /popup Main /Just L /Text Koordi�   natensysteme!�E /L /Jump Objekte /Link /Macro /Play /popup �   Main /Just L /Text Objekte!�Q /L /Jump Objektklassen /Link �   /Macro /Play /popup Main /Just L /Text Objektklassen!�� /L �   /Jump Selektierte und aktivierte Objekte /Link /Macro /Play    /popup Main /Just L /Text Recherchierte, selektierte und a  ktivierte Objekte!� /P /Just L /Text ��!� /H /Just L /Tex  te!� /P /Just L /Text !�] /L /Jump Was ist ein Objekt /Lin�  t Reference!�G /L /Jump Anhang A /Link /Macro /Play /popup    gespeicherten raumbezogenen und sachbezogenen Daten. Gleic  hzeitig kann es �ber thematische Relationen in Verbindung m  it anderen Objekten stehen.����Grunds�tzlich werden untersc�   hieden:!� /B /Just L /Text Punktobjekt!� /B /Just L /Text  bjekt;Fl�chenobjekt;Linienobjekt;Punktobjekt;�� N�     �	  .  G�� 
Q  * 1 J     � Topic@Objekte  �    �  
  	  � 1010   �  ��8Y     �  �� Cp     � Objekte��   R�     �  �� 	b%  � -�   !� /T N /Just L /Text Objek$  eine vorgebbare Fl�chensignatur.!�. Fl�chensignatur,(Global  seln'). Die Darstellung eines Fl�chenobjektes erfolgt �ber �   �  �^�� 
|  5 < U     � Topic@Was ist ein Objekt %   Was ist ein Objekt�� ]�     �  �� 	�y  �-�   !�' /     ?  
y �                                                   k /Macro /Play /popup Main /Just L /Text Was ist ein Objekt6   emnach die M�glichkeit der gleichzeitigen Analyse seiner La!    �  �� �     �  ��>[     �  �� Ex     � Punktsig  �   ��� 
@  0 7 L     � Topic@Punktsignatur  �  /   dessen Raumbezug in Form eines zu einer Fl�che geschlossen  ekt,(Global), 0,Ein Fl�chenobjekt ist ein Objekt in TRiAS�,  lobjekte.!�  Datenimport,(Global), 0,<(None)>!�QFl�chenobj  stellten Darstellungsparametern der Objektklassen und Einze  ener Objektklassen im TRiAS�-Fenster entsprechend den einge  .!�� Ansicht,(Global), 2,Darstellung aller Objekte vorgegeb  also blinkt und durch ein Fokus-Rechteck gekennzeichnet ist  ist und dort das vom Nutzer derzeit aktivierte Objekt ist,   einer Operation in einem Objekt-Recherchefenster enthalten     bjekten.  
� �                                             ��Ein Objekt in TRiAS� repr�sentiert die Einheit der zu ein  em in der realen Welt existierenden Vorgang oder Gegenstand  ge, seiner Eigenschaften und seiner Verbindung zu anderen O0  natur�� T�     �  �� 	d�   * -�   !�  /T N /Just L /Te1  text f�r einen Identifikator, ein Merkmal oder eine Relatio"  st ein Identifikator>!�� Kurztext,(Global), 2,Beschreibungs#  ), 2,<Flaechensignatur>!�5 Identifikator,(Global), 2,<Was i  T N /Just L /Text Was ist ein Objekt ?!�?/P /Just L /Text      /Text Fl�chensignatur  
� �  � 1003                   &  hensignatur�� W�     �  �� 	g�   * -�   !�  /T /Just L'      �  �� �     �  ��A^     �  �� H~     � Flaec(  �   ���� 
E  3 : O     � Topic@Flaechensignatur  �+  �   �`�� 
�  1 8 Q     � Topic@Liniensignatur  �  ,    �  	  � 1009   �  ��?`     �  �� J~     � Lin-  iensignatur�� Y�     �  �� 	i�   ) -�   !� /T /Just L     /Text Liniensignatur  
� �                                 Polygonzug weitere zugeh�rige Polygone enthalten kann ('In.  en Polygonzuges (Punktfolge) dargestellt wird, wobei dieser    xt Punktsignatur  
� �  � 1012                         n@  n, der maximal 32 Zeichen umfassen kann und im allgemeinen A  Identifikator /Link /Macro /Play /popup Main /Just L /Text 2   /Text Was ist eine Objektklasse ?!�k /L /Jump Was ist ein 3  st eine Objektklasse /Link /Macro /Play /popup Main /Just LL  tifikator!�c/P /Just L /Text Der Unterschied zwischen dem 5  1 /Just L /Text Unterschiede zwischen Objektklasse und Iden6  rgabe seiner grundlegenden Darstellungsparameter. ��!�G /S 7  ist wichtig f�r seine Zuordnung zu einer Ansicht und zur Vo[  doch die Lesbarkeit  z.B. der Legende.����Prinzipiell k�nne9  reibungstext (Langtext) mu� nicht definiert sein, erh�ht je:  nsdarstellung und mu� daher definiert sein. Der lange Besch;  et. Er dient einer schnellen und �bersichtlichen Informatio<  t (Kurztext) wird in den meisten Dialogen in TRiAS� verwendK  ator, ein Merkmal oder eine Relation, der beliebig viele Ze>  bal), 2,Ausf�hrlicher Beschreibungstext f�r einen Identifik?  eine schlagwortartige Bezeichnung enth�lt.!�� Langtext,(Glo    Was ist ein Identifikator ?  
� �                        C  �Jedem dieser Schl�ssel kann ein kurzer und ein langer Besc=  hreibungstext zugeordnet werden. Der kurze Beschreibungstex\  nsignatur>!�' Objekt,(Global), 2,<Was ist ein Objekt>!�9 ObD  ebbare Liniensignatur.!�+ Liniensignatur,(Global), 2,<LinieE  Die Darstellung eines Linienobjektes erfolgt �ber eine vorgF  ines einzelnen Polygonzuges (Punktfolge) dargestellt wird. G  objekt ist ein Objekt in TRiAS�, dessen Raumbezug in Form eH  zeichnung enth�lt.
!�� Linienobjekt,(Global), 2,Ein Linien�   /P /Just L /Text ��Eine Objektklasse ist eine logische ZusI  ichen umfassen kann und im allgemeinen eine vollst�ndige Beo  Begriff 'Objektklasse' und dem Begriff Identifikator' besteJ  2-�   !�, /T N /Just L /Text Was ist eine Objektklasse!�FM      � Was ist eine Objektklasse�� d�     �  �� 	t�  N  asse  �    �  	  � 1017   �  ��Jk     �  �� U� O  �  y�� 
y  < C \   $  � Topic@Was ist eine Objektkl�B  d z.B. "Wald", "Stra�e", "Flu�", "Betriebsgel�nde" etc.)���S  �,/P /Just L /Text ��Um gro�e Mengen von Objekten handhabbT  ar verwalten zu k�nnen, wird in TRiAS� jedem Objekt ein Ide]  ntifikator zugeordnet. Dieser Identifikator ist ein 8-10 stp  tenform einige Informationen �ber eine Menge von Objekten eU  ektrecherchefenster,(Global), 2,Ein Fenster, welches in LisV  Objektklasse,(Global), 2,<Was ist eine Objektklasse>!�� Obj    m Potsdam  
� �                                          X   die Verwendung der durch die uve GmbH FernerkundungszentruY  ation der Objekte verwendet werden. Es empfielt sich jedochZ   beliebige Zahlenschl�ssel zur Identifikation und KlassifikW  jekte,Was ist eine Objektklasse, 0,<Was ist ein Objekt>!�4 ^  elliger hierarchischer Zahlenschl�ssel, der in �bereinstimm_  ung mit dem zentralen Merkmal eines Objektes vergeben wird.`    Er wird h�ufig zur Zuordnung von Objekten zu einer thematQ  ischen Objektklasse verwendet (typische Identifikatoren sinm   'Wald' oder 'Stra�e' zu sein) ist, eine Objektklasse dagegq  -Recherchefenster enthalten ist und dort vom Nutzer ausgew�b   2,Ein Objekt, welches nach einer Operation in einem Objektc   Lage zu anderen Objekten.!�� selektiertes Objekt,(Global),d  zug,(Global), 2,Die Form und Gr��e eines Objektes sowie diee  tur.!�) Punktsignatur,(Global), 2,<Punktsignatur>!�[ Raumbef  eines Punktobjektes erfolgt �ber eine vorgebbare Punktsignag   eines einzelnen Punktes dargestellt wird. Die Darstellung h  ktobjekt ist ein Objekt in TRiAS�, dessen Raumbezug in Formi  e zusammengestellt wird.!�� Punktobjekt,(Global), 2,Ein Pun�  al ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�;  ,    ien sein kann.  
� �                                     l  en eine Zusammenfassung von Objekten nach beliebigen Kritera   Klassifikation von Objekte nach deren Hauptmerkmal  (z.B.:n  ht darin, da� ein Identifikator ein Zahlenschl�ssel f�r diej  nth�lt, die im Ergebnis eines Kommandos oder einer RecherchB�  hlt wurde (in der Listbox gekennzeichnet also selektiert iss    L-�   !�- /T N /Just L /Text Koordinaten der Datenbasis�  !�H/P /Just L /Text ��Die Koordinaten der Objekte, die in u   N /Just L /Text Inhaltsverzeichnis!�" /H /Just L /Text All�   gemeine Fragen!�s /L /Jump Darstellung /Link /Macro /Play /w  �  z�� 
�  5 < U     � Topic@Koordinatensysteme x   �    �  	  � 1008   �  ��Cd     �  �� N�     �y   Koordinatensysteme�� ]�     �  �� 	m�  -�   !�% /Tz   N /Just L /Text Koordinatensysteme!� /P /Just L /Text !�k{   /L /Jump Koordinaten der Datenbasis /Link /Macro /Play /po|  pup Main /Just L /Text Koordinaten der Datenbasis!�c /L /Ju�  mp Angezeigte Koordinaten /Link /Macro /Play /popup Main /J~     a��� 
~  < C \   $  � Topic@Was ist ein Identifik  ator  �    �  	  � 1015   �  ��Jk     �  �� U� �      � Was ist ein Identifikator�� d�     �  �� 	t  R  h-�   !�. /T N /Just L /Text Was ist ein Identifikator ?!r       � Koordinaten der Datenbasis�� e�     �  �� 	u��  m Koordinatensystem keine Sprunghaften Ver�nderungen der Ko�  tetig bedeutet, da� bei einer ebenm��igen Lagever�nderung i�  t, welches stetig und orthogonal ist.!�� /B /Just L /Text S�  e Objektgeometrien immer in einem Koordinatensystem abgeleg�   einfache Verwaltung der Koordinaten zu erm�glichen sind di�   immer den angezeigten Koordinaten.����Um eine homogene und�  der TRiAS�-Datenbasis abgespeichert sind, entsprechen nicht�  _  0}�� 
�  9 @ Y   !  � Topic@Angezeigte Koordinate    ust L /Text Angezeigte Koordinaten  
� �                 �    {k�� 
�  = D ]   %  �  Topic@Koordinaten der Daten�   L /Text ��Die angezeigten bzw. bei einer Eingabe erwartete�   !�) /T N /Just L /Text Angezeigte Koordinaten!�v /P /Just�    � Angezeigte Koordinaten�� a�     �  �� 	qV  � -�  �  n  �    �  	  � 1000   �  ��Gh     �  �� R�   �  basis  �    �  	  � 1007   �  ��Kl     �  �� V�n�  ordinatenwerte auftreten. Da� ist beispielsweise bei einem �  ojekt unter dem angegebenen Namen und wird sofort wieder an�  as Hauptfenster angezeigt wird, erzeugt ein neues TRiAS�-Pr�  ame!�� /P 1 /Just L /Text TRiAS� wird gestartet, ohne da� d�  \NAME\NAME.RIS' gesucht.!�" /B 1 /Just L /Text /init Datein                                                               �  n Koordinaten sind (in gewissen Grenzen) vorgebbar.  
� �    e den bereits erfassten Daten entsprechen.  
� �         �  r Daten aus Korrdinatensystemen verwendet werden d�rfen, di�  chten, da� bei zus�tzlicher Datenerfassung (Datenimport) nu�  Umrechnung vorgenommen. Ferner ist es jedoch wichtig zu bea�  ge bzw. bei der Eingabe von Koordinaten eine entsprechende �   L /Text Um diesen Kriterien zu gen�gend wird bei der Anzei�  chsen des Systemes senkrecht aufeinanderstehen.!�Y/P /Just�   /B /Just L /Text Orthogonal bedeutet, da� die Koordinatena�  Streifenwechsel in allen Gau�-/Kr�ger-Systemen der Fall.!�it   Inhaltsverzeichnis�� ]�     �  �� 	m�  D-�   !�% /T�   /Text Der angegebene Dateiname wird als Projektname verwen�  det, und TRiAS� versucht dieses Projekt sofort zu er�ffnen.�  !�v/P 2 /Just L /Text Ist kein vollst�ndiger Pfad gegeben,�   so wird das Projekt in einem Unterverzeichnis des Standard�  - Projektverzeichnisses gesucht, welches den Namen des Proj�  ektes tr�gt.��z.B. Bei einem Standard- Projektverzeichnis '�  1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  �   Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !��  C:\TRIAS\PROJEKTE' und einem angegebenen Dateinamen 'NAME.R�  IS', so wird das Projekt unter dem Namen 'C:\TRIAS\PROJEKTE�  tfenster angezeigt wird, zeigt ein Dialogfenster an, in dem�  /P 1 /Just L /Text TRiAS� wird gestartet, ohne da� das Haup�  hen Vorgaben, wie oben.!� /B 1 /Just L /Text /init:ask!�� �  gehalten. Bei fehlemdem vollst�ndigen Pfad gelten die gleic�   ein Projektname direkt vorgegeben werden kann. Dieses TRiAB�  ben werden:!� /B 1 /Just L /Text Dateiname!�� /P 1 /Just L�   Dateinamen sinnvoll)!�N /P 1 /Just L /Text Das gegebene TR�  rtfenster angezeigt wird!�4 /B 1 /Just L /Text /r �(nur mit�  Just L /Text TRiAS� wird gestartet, jedoch ohne da� das Sta�  ofort wieder angehalten.!� /B 1 /Just L /Text /n!�Y /P 1 /�  -Projekt mit dem gegebenen Namen auf dem Desktop und wird s�  � das Hauptfenster angezeigt wird, erzeugt ein neues TRiAS��  ows95)!�� /P 1 /Just L /Text TRiAS� wird gestartet, ohne da�  n.!�; /B 1 /Just L /Text /init:desktop Dateiname �(nur Wind�  S�-Projekt wird erzeugt, anschlie�end wird TRiAS� angehalte�  v
  ���� 
�  9 @ Y   !  � Topic@Komandozeilenparamete�  r  �    �  	  � 1006   �  ��Gh     �  �� R�   �    � Komandozeilenparameter�� a�     �  �� 	qm
  �	-�  �   !�) /T N /Just L /Text Komandozeilenparameter!�N /P /Just    ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�            �   L /Text ��Es k�nnen folgende Komandozeilenparameter angege�  iAS�-Projekt wird schreibgesch�tzt er�ffnet.!� /B 1 /Just �    �    �  	  � 1002   �  ��De     �  �� O�     ��  �  �y�� 
�  6 = V     � Topic@Doppelte Menupunkte    �scht werden soll.  
� �                                 �  n sollte benutzt werden, bevor TRiAS� von einem rechner gel�  ren. Anschlie�end wird das Programm angehalten. Diese Optio�  die f�r die w�hrend der Arbeit mit dem Programmnotwendig wa�  estartet und bereinigt alle eingerichteten Systemeintr�ge, �  st L /Text /unregserver!�/P 1 /Just L /Text TRiAS� wird g�  ebene Standardansicht wird nicht initialisiert.!� /B 1 /Ju�  t Das gegebene TRiAS�-Projekt wird er�ffnet. Eine evtl. geg�  /Text /s�(nur mit Dateinamen sinnvoll)!�{ /P 1 /Just L /Tex�  Anschlie�end wird das Programm angehalten.!�3 /B 1 /Just L �  r die richtige Funktion des Programmes notwendig sind ein. �  tet und richtet alle notwendigen Systemeintr�ge ein, die f��  L /Text /regserver!�� /P 1 /Just L /Text TRiAS� wird gestar�   Doppelte Menupunkte�� ^�     �  �� 	n�  	-�   !�( �  e und aktivierte Objekte!�/P /Just L /Text ��Im Resultat �      �  �� 	}  K-�   !�5 /T N /Just L /Text Selektiert�   �� ^�   '  �" Selektierte und aktivierte Objekte�� m� �  �  &��� 
�  5 < U     � Topic@Inhaltsverzeichnis �   �    �  	  � 1005   �  ��Cd     �  �� N�     ��  erten Objekte dieses Fensters, je nach dem, ob das ausgew�h�  ch entweder auf das aktivierte Objekt oder auf alle selekti�  �Menupunkte im Menu des Objektrecherchefensters beziehen si�  er aktuellen Ansicht und des aktuellen Bildausschnittes.����  uf eine  oder mehrere Objektklassen oder auf alle Objekte d�  beziehen sich die Menupunkte/Kommandos im Hauptmenu immer a�  h im Menu aller Objektrecherchefenster enthalten.����Dabei �  e der Menupunkte/Kommandos sind sowohl im Hauptmenu als auc�  t ��Warum gibt es in TRiAS� 'doppelte Menupunkte' ?����Viel�  /T N /Just L /Text Doppelte Menupunkte ?!�%/P /Just L /Texn�  einer Recherche oder anderweitigen Operation kann ein Objek�    ���� 
�  E L e   -  �( Topic@Selektierte und aktiv�  ierte Objekte  �    �  	  � 1013   �  ��St     �       !�  !�  !�                                               �   !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !��  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !� �  kte k�nnen mit beliebigen Fonts dargestellt werden.!�  !�  �  ls zus�tzliche Signatur anderer Objekte in TRiAS�. Textobje�  ealen Welt hat. Es dient der textlichen Beschreibung oder a�   in TRiAS�, welches im allgemeinen kein �quivalent in der r�  t..!�Textobjekt,(Global), 0,Ein Textobjekt ist ein Objekt�  te' bezeichnet.����Nach Erzeugen dieses Fensters ist genau �  Fenster enthaltenen Objekte werden als 'recherchierte Objek�  trecherchefenster erzeugt werden. Alle in einem derartigen   /Play /popup Main /Just L /Text Index!�_ /L /Jump Stichwort�  Main /Just L /Text Anhang A!�A /L /Jump Index /Link /Macro n   lte Kommando sich von seinem Inhalt her auf ein oder mehrer  en mit der rechten Maustaste lassen sich in diesem Objektre�  iges Bet�tigen der Control-Taste (Strg bzw. Ctrl) und Klick�  eichzeitig auch aktiviert ist (blinkt).����Durch gleichzeit�  ein Objekt 'selektiert' (unterlegt), wobei dieses Objekt gl    nstellungen f�r den betreffenden Dialog.  
� �           �  alisierung, das aktivierte Objekt dagegen liefert die Vorei�  c.) erhalten alle selektierten Objekte die ausgew�hlte Visu�  isualisierung (Darstellungsparameter wie Farbe, Signatur et�  �/B /Just L /Text Beim Einstellen einer objektbezogenen V�  n die selektierten Objekte immer die geschnittenenen sind.!�  chnitt das aktivierte Objekte immer das schneidende, wogege�   Hier einige Beispiele:!�� /B /Just L /Text Beim Objektvers�  pielt das aktivierte Objekt die Rolle eines Bezugsobjektes.�  gew�hlte Menupunkt auf alle selektierten Objekte bezieht, s�  e Objekte bezieht.����Selbst dann jedoch, wenn sich des ausB  cherchefenster unabh�ngig voneinander einzelne Objekte sele  isualiserungsfehler�� [�     �  �� 	k\  � -�   !�' /T   N /Just L /Text Visualiserungsfehler!�� /P /Just L /Text W  arum werden fehlende Visualiserungen nicht gemeldet, obwohl   das 'H�kchen' f�r das Ignorieren wieder entfernt wurde ?      
� �                                                         ichwortverzeichnis  
� �                                   verzeichnis /Link /Macro /Play /popup Main /Just L /Text St
  g�� R�     �  �� 	bl  � -�   !�+ /T N /Just L /Text D  arstellung von Objekten!�@ /H /Just L /Text Farbe, Signatur  en, Darstellungsreihenfolge etc.!�` /L /Jump Visualiserungs  fehler /Link /Macro /Play /popup Main /Just L /Text Visuali    nze Bereiche von Objekte selektieren.  
� �                s Bet�tigen der Shift-Taste (Umschalt-Taste) lassen sich ga  ckte Objekt aktiviert wird (blinkt).����Durch gleichzeitige  ktieren (unterlegen), wobei nur das jeweils zuletzt angekli    �    �    �    �  ��Eb     �  �� L�     � V                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     sierungsfehler  
} �                                       u  �2�� 
�  . 5 J     � Topic@Darstellung  �   	   �    �    �  ��<Y     �  �� Ct     � Darstellun  e  �S�� 
�  7 > S     � Topic@Visualiserungsfehler